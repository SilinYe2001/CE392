

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO key_generation 
  PIN clk 
    ANTENNAPARTIALMETALAREA 1.0976 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6256 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 32.0513 LAYER metal4 ; 
    ANTENNAMAXAREACAR 55.1275 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 221.461 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 1.12129 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAGATEAREA 32.0513 LAYER metal5 ; 
    ANTENNAMAXAREACAR 55.1282 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 221.466 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.1219 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 1.7052 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER metal6 ;
    ANTENNAGATEAREA 32.0775 LAYER metal6 ; 
    ANTENNAMAXAREACAR 55.1813 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 221.681 LAYER metal6 ;
    ANTENNAMAXCUTCAR 2.05333 LAYER via6 ;
  END clk
  PIN rst 
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.294 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 18.3848 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 73.8528 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.29925 LAYER metal6 ; 
    ANTENNAMAXAREACAR 196.329 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 792.002 LAYER metal6 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via6 ;
  END rst
  PIN start 
    ANTENNAPARTIALMETALAREA 0.6468 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6656 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.3908 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.6416 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 26.5776 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 106.467 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 555.847 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 2230.14 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END start
  PIN p[63] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.55375 LAYER metal7 ; 
    ANTENNAMAXAREACAR 30.3723 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 121.574 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.03709 LAYER via7 ;
  END p[63]
  PIN p[62] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.45675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 35.3328 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 141.806 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.03956 LAYER via7 ;
  END p[62]
  PIN p[61] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 52.1858 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 211.042 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.79431 LAYER via7 ;
  END p[61]
  PIN p[60] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 146.228 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 588.575 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41963 LAYER via7 ;
  END p[60]
  PIN p[59] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.464 LAYER metal7 ; 
    ANTENNAMAXAREACAR 158.155 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 636.438 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.17033 LAYER via7 ;
  END p[59]
  PIN p[58] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 63.8141 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 258.256 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.13829 LAYER via7 ;
  END p[58]
  PIN p[57] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.464 LAYER metal7 ; 
    ANTENNAMAXAREACAR 90.1521 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 364.101 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.42009 LAYER via7 ;
  END p[57]
  PIN p[56] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.255 LAYER metal7 ; 
    ANTENNAMAXAREACAR 77.4061 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 313.373 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.42232 LAYER via7 ;
  END p[56]
  PIN p[55] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.673 LAYER metal7 ; 
    ANTENNAMAXAREACAR 40.0179 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 163.821 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41841 LAYER via7 ;
  END p[55]
  PIN p[54] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.30725 LAYER metal7 ; 
    ANTENNAMAXAREACAR 70.7704 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 286.597 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.79681 LAYER via7 ;
  END p[54]
  PIN p[53] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.30725 LAYER metal7 ; 
    ANTENNAMAXAREACAR 72.059 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 291.97 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.42169 LAYER via7 ;
  END p[53]
  PIN p[52] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 104.494 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 421.661 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.79474 LAYER via7 ;
  END p[52]
  PIN p[51] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 71.2419 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 286.3 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41963 LAYER via7 ;
  END p[51]
  PIN p[50] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 54.0096 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 218.119 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04451 LAYER via7 ;
  END p[50]
  PIN p[49] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.647 LAYER metal7 ; 
    ANTENNAMAXAREACAR 110.44 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 445.106 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.4186 LAYER via7 ;
  END p[49]
  PIN p[48] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 103.816 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 418.73 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41963 LAYER via7 ;
  END p[48]
  PIN p[47] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 108.577 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 437.689 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.79474 LAYER via7 ;
  END p[47]
  PIN p[46] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 55.3823 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 223.703 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04407 LAYER via7 ;
  END p[46]
  PIN p[45] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.647 LAYER metal7 ; 
    ANTENNAMAXAREACAR 64.2099 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 260.189 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.8875 LAYER via7 ;
  END p[45]
  PIN p[44] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.41175 LAYER metal7 ; 
    ANTENNAMAXAREACAR 40.9424 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 166.284 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.42058 LAYER via7 ;
  END p[44]
  PIN p[43] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 39.3207 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 160.789 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41919 LAYER via7 ;
  END p[43]
  PIN p[42] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 46.2521 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 191.683 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.88809 LAYER via7 ;
  END p[42]
  PIN p[41] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 60.5922 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 246.053 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41963 LAYER via7 ;
  END p[41]
  PIN p[40] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 32.0704 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 131.55 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04407 LAYER via7 ;
  END p[40]
  PIN p[39] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.464 LAYER metal7 ; 
    ANTENNAMAXAREACAR 41.1276 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 165.66 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04497 LAYER via7 ;
  END p[39]
  PIN p[38] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 46.1352 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 187.877 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04407 LAYER via7 ;
  END p[38]
  PIN p[37] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.69925 LAYER metal7 ; 
    ANTENNAMAXAREACAR 47.9164 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 195.145 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41823 LAYER via7 ;
  END p[37]
  PIN p[36] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.464 LAYER metal7 ; 
    ANTENNAMAXAREACAR 48.3837 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 197.177 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04497 LAYER via7 ;
  END p[36]
  PIN p[35] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 37.8974 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 153.255 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.819434 LAYER via7 ;
  END p[35]
  PIN p[34] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.62075 LAYER metal7 ; 
    ANTENNAMAXAREACAR 32.1815 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 129.304 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.527883 LAYER via7 ;
  END p[34]
  PIN p[33] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5425 LAYER metal7 ; 
    ANTENNAMAXAREACAR 47.2204 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 191.136 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.910314 LAYER via7 ;
  END p[33]
  PIN p[32] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 32.5803 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 132.041 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.856946 LAYER via7 ;
  END p[32]
  PIN p[31] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.72525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 20.0759 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 80.6209 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.442293 LAYER via7 ;
  END p[31]
  PIN p[30] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 25.8766 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 105.507 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.903405 LAYER via7 ;
  END p[30]
  PIN p[29] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 24.2101 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 97.8558 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.559951 LAYER via7 ;
  END p[29]
  PIN p[28] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.647 LAYER metal7 ; 
    ANTENNAMAXAREACAR 35.3016 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 141.472 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.730681 LAYER via7 ;
  END p[28]
  PIN p[27] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 125.63 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 506.095 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41919 LAYER via7 ;
  END p[27]
  PIN p[26] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 19.9531 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 80.9844 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.535085 LAYER via7 ;
  END p[26]
  PIN p[25] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 23.2363 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 94.3937 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.697811 LAYER via7 ;
  END p[25]
  PIN p[24] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 75.1814 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 304.41 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41963 LAYER via7 ;
  END p[24]
  PIN p[23] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 18.8958 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 75.9814 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.619793 LAYER via7 ;
  END p[23]
  PIN p[22] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7515 LAYER metal7 ; 
    ANTENNAMAXAREACAR 34.3657 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 138.744 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.73017 LAYER via7 ;
  END p[22]
  PIN p[21] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 33.0677 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 134.351 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.794426 LAYER via7 ;
  END p[21]
  PIN p[20] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.464 LAYER metal7 ; 
    ANTENNAMAXAREACAR 20.843 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 84.1205 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.13875 LAYER via7 ;
  END p[20]
  PIN p[19] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 20.4547 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 82.8301 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.688698 LAYER via7 ;
  END p[19]
  PIN p[18] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.647 LAYER metal7 ; 
    ANTENNAMAXAREACAR 66.297 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 266.619 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.79372 LAYER via7 ;
  END p[18]
  PIN p[17] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.41175 LAYER metal7 ; 
    ANTENNAMAXAREACAR 51.6128 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 207.284 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04546 LAYER via7 ;
  END p[17]
  PIN p[16] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 83.2569 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 336.587 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41963 LAYER via7 ;
  END p[16]
  PIN p[15] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 65.661 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 266.425 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.32541 LAYER via7 ;
  END p[15]
  PIN p[14] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 129.916 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 523.192 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41963 LAYER via7 ;
  END p[14]
  PIN p[13] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.41175 LAYER metal7 ; 
    ANTENNAMAXAREACAR 56.4343 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 228.688 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.13924 LAYER via7 ;
  END p[13]
  PIN p[12] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 31.6617 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 127.098 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04451 LAYER via7 ;
  END p[12]
  PIN p[11] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.62075 LAYER metal7 ; 
    ANTENNAMAXAREACAR 32.3839 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 131.495 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04367 LAYER via7 ;
  END p[11]
  PIN p[10] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 76.3056 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 307.27 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41963 LAYER via7 ;
  END p[10]
  PIN p[9] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.51625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 59.1018 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 237.003 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.950726 LAYER via7 ;
  END p[9]
  PIN p[8] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.464 LAYER metal7 ; 
    ANTENNAMAXAREACAR 91.1729 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 366.239 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04497 LAYER via7 ;
  END p[8]
  PIN p[7] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5685 LAYER metal7 ; 
    ANTENNAMAXAREACAR 57.1958 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 230.333 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04407 LAYER via7 ;
  END p[7]
  PIN p[6] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.41175 LAYER metal7 ; 
    ANTENNAMAXAREACAR 42.1067 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 172.023 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04546 LAYER via7 ;
  END p[6]
  PIN p[5] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3595 LAYER metal7 ; 
    ANTENNAMAXAREACAR 43.0656 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 174.264 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.42112 LAYER via7 ;
  END p[5]
  PIN p[4] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.59475 LAYER metal7 ; 
    ANTENNAMAXAREACAR 50.6484 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 203.778 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.41899 LAYER via7 ;
  END p[4]
  PIN p[3] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.59475 LAYER metal7 ; 
    ANTENNAMAXAREACAR 42.2352 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 170.849 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04387 LAYER via7 ;
  END p[3]
  PIN p[2] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.38575 LAYER metal7 ; 
    ANTENNAMAXAREACAR 31.0271 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 124.857 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04572 LAYER via7 ;
  END p[2]
  PIN p[1] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.27375 LAYER metal7 ; 
    ANTENNAMAXAREACAR 59.6001 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 240.381 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.32154 LAYER via7 ;
  END p[1]
  PIN p[0] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.73625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 95.4051 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 385.849 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.47854 LAYER via7 ;
  END p[0]
  PIN q[63] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2355 LAYER metal7 ; 
    ANTENNAMAXAREACAR 105.69 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 425.286 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.784898 LAYER via7 ;
  END q[63]
  PIN q[62] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.4165 LAYER metal7 ; 
    ANTENNAMAXAREACAR 25.7873 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 105.085 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.939924 LAYER via7 ;
  END q[62]
  PIN q[61] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 29.8388 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 122.104 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.76994 LAYER via7 ;
  END q[61]
  PIN q[60] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 78.2859 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 314.766 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.578397 LAYER via7 ;
  END q[60]
  PIN q[59] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.44275 LAYER metal7 ; 
    ANTENNAMAXAREACAR 16.698 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 68.9701 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690225 LAYER via7 ;
  END q[59]
  PIN q[58] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 31.8426 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 129.081 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.01962 LAYER via7 ;
  END q[58]
  PIN q[57] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 72.9212 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 294.257 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.989858 LAYER via7 ;
  END q[57]
  PIN q[56] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.49475 LAYER metal7 ; 
    ANTENNAMAXAREACAR 38.1961 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 154.976 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.939873 LAYER via7 ;
  END q[56]
  PIN q[55] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 60.673 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 245.783 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.01962 LAYER via7 ;
  END q[55]
  PIN q[54] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 85.3037 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 343.423 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.989858 LAYER via7 ;
  END q[54]
  PIN q[53] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 18.2544 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 73.1772 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.534123 LAYER via7 ;
  END q[53]
  PIN q[52] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 65.7244 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 265.989 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.01962 LAYER via7 ;
  END q[52]
  PIN q[51] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 79.1372 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 319.39 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.989858 LAYER via7 ;
  END q[51]
  PIN q[50] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 20.4489 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 83.2093 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690174 LAYER via7 ;
  END q[50]
  PIN q[49] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 66.2939 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 267.934 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.01962 LAYER via7 ;
  END q[49]
  PIN q[48] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 63.7861 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 257.717 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.740176 LAYER via7 ;
  END q[48]
  PIN q[47] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.495 LAYER metal7 ; 
    ANTENNAMAXAREACAR 14.4644 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 58.1348 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690191 LAYER via7 ;
  END q[47]
  PIN q[46] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 71.5412 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 288.923 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.01962 LAYER via7 ;
  END q[46]
  PIN q[45] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 84.1513 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 339.392 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.989858 LAYER via7 ;
  END q[45]
  PIN q[44] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.495 LAYER metal7 ; 
    ANTENNAMAXAREACAR 18.201 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 73.3549 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690191 LAYER via7 ;
  END q[44]
  PIN q[43] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 39.9028 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 160.558 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.552115 LAYER via7 ;
  END q[43]
  PIN q[42] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 58.0037 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 233.657 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.615873 LAYER via7 ;
  END q[42]
  PIN q[41] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 18.732 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 75.7184 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690174 LAYER via7 ;
  END q[41]
  PIN q[40] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 82.1361 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 331.302 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.01962 LAYER via7 ;
  END q[40]
  PIN q[39] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 119.881 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 482.097 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.989858 LAYER via7 ;
  END q[39]
  PIN q[38] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 17.4258 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 70.1066 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690174 LAYER via7 ;
  END q[38]
  PIN q[37] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 38.0238 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 153.423 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.552115 LAYER via7 ;
  END q[37]
  PIN q[36] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 40.1014 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 162.82 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.578397 LAYER via7 ;
  END q[36]
  PIN q[35] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 18.6322 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 75.2932 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.03513 LAYER via7 ;
  END q[35]
  PIN q[34] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 33.4361 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 134.463 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.520856 LAYER via7 ;
  END q[34]
  PIN q[33] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 50.9212 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 205.41 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.616032 LAYER via7 ;
  END q[33]
  PIN q[32] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 23.8193 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 94.7128 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.431929 LAYER via7 ;
  END q[32]
  PIN q[31] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 36.3911 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 147.232 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.552115 LAYER via7 ;
  END q[31]
  PIN q[30] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 52.2869 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 210.33 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.605667 LAYER via7 ;
  END q[30]
  PIN q[29] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.57325 LAYER metal7 ; 
    ANTENNAMAXAREACAR 16.9705 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 68.1491 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690141 LAYER via7 ;
  END q[29]
  PIN q[28] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 17.2573 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 70.6631 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.739675 LAYER via7 ;
  END q[28]
  PIN q[27] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 25.7093 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 104.823 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.672177 LAYER via7 ;
  END q[27]
  PIN q[26] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 13.3634 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 54.8134 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690174 LAYER via7 ;
  END q[26]
  PIN q[25] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 23.2514 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 94.3581 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.552115 LAYER via7 ;
  END q[25]
  PIN q[24] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 32.2815 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 130.814 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.605667 LAYER via7 ;
  END q[24]
  PIN q[23] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 18.0609 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 72.8775 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.471703 LAYER via7 ;
  END q[23]
  PIN q[22] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 47.0482 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 189.537 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.552115 LAYER via7 ;
  END q[22]
  PIN q[21] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 41.6033 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 168.474 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.709812 LAYER via7 ;
  END q[21]
  PIN q[20] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 17.9547 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 72.4905 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.939856 LAYER via7 ;
  END q[20]
  PIN q[19] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 52.0125 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 209.142 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.458336 LAYER via7 ;
  END q[19]
  PIN q[18] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 36.6562 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 146.863 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.535711 LAYER via7 ;
  END q[18]
  PIN q[17] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.57325 LAYER metal7 ; 
    ANTENNAMAXAREACAR 13.7616 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 55.0044 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690141 LAYER via7 ;
  END q[17]
  PIN q[16] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 21.0514 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 85.7062 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.552115 LAYER via7 ;
  END q[16]
  PIN q[15] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 23.1061 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 93.4074 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.549163 LAYER via7 ;
  END q[15]
  PIN q[14] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.495 LAYER metal7 ; 
    ANTENNAMAXAREACAR 22.762 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 90.3546 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690191 LAYER via7 ;
  END q[14]
  PIN q[13] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 33.0021 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 133.59 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.552115 LAYER via7 ;
  END q[13]
  PIN q[12] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 27.9409 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 112.624 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.361604 LAYER via7 ;
  END q[12]
  PIN q[11] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.521 LAYER metal7 ; 
    ANTENNAMAXAREACAR 14.8864 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 59.6446 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.690174 LAYER via7 ;
  END q[11]
  PIN q[10] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 24.8184 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 100.725 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.458336 LAYER via7 ;
  END q[10]
  PIN q[9] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 30.9162 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 124.901 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.455383 LAYER via7 ;
  END q[9]
  PIN q[8] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.57325 LAYER metal7 ; 
    ANTENNAMAXAREACAR 16.0971 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 64.6933 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.461266 LAYER via7 ;
  END q[8]
  PIN q[7] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ; 
    ANTENNAMAXAREACAR 39.1501 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 158.385 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.458336 LAYER via7 ;
  END q[7]
  PIN q[6] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 35.4751 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 142.983 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.455383 LAYER via7 ;
  END q[6]
  PIN q[5] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.75275 LAYER metal7 ; 
    ANTENNAMAXAREACAR 19.914 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 80.1611 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.04276 LAYER via7 ;
  END q[5]
  PIN q[4] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 39.4057 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 159.243 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.361604 LAYER via7 ;
  END q[4]
  PIN q[3] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.366 LAYER metal7 ; 
    ANTENNAMAXAREACAR 25.9172 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 105.091 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.361604 LAYER via7 ;
  END q[3]
  PIN q[2] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.57075 LAYER metal7 ; 
    ANTENNAMAXAREACAR 58.645 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 235.274 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.537931 LAYER via7 ;
  END q[2]
  PIN q[1] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.28775 LAYER metal7 ; 
    ANTENNAMAXAREACAR 100.139 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 402.671 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.932535 LAYER via7 ;
  END q[1]
  PIN q[0] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.39225 LAYER metal7 ; 
    ANTENNAMAXAREACAR 111.665 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 448.41 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.668413 LAYER via7 ;
  END q[0]
  PIN done 
    ANTENNAPARTIALMETALAREA 0.3332 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4112 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.3916 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6448 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 22.5596 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 90.3168 LAYER metal6 ;
  END done
  PIN mem_wr_en 
    ANTENNAPARTIALMETALAREA 0.0399 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1596 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2548 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0976 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.7428 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0496 LAYER metal6 ;
  END mem_wr_en
  PIN addr_rd_out[63] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.4777 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9304 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.13075 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.2871 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 69.1428 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[63]
  PIN addr_rd_out[62] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.0752 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.6699 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 42.8261 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[62]
  PIN addr_rd_out[61] 
    ANTENNAPARTIALMETALAREA 0.0798 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3192 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal4 ; 
    ANTENNAMAXAREACAR 11.7323 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 47.0793 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via4 ;
  END addr_rd_out[61]
  PIN addr_rd_out[60] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.6097 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4388 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.94542 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 38.6208 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[60]
  PIN addr_rd_out[59] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5628 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2708 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.83659 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 38.1128 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[59]
  PIN addr_rd_out[58] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.6125 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4696 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.82399 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 38.0475 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.24998 LAYER via3 ;
  END addr_rd_out[58]
  PIN addr_rd_out[57] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5327 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1504 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.4571 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 52.8451 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[57]
  PIN addr_rd_out[56] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.61355 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4934 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.7616 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.2605 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[56]
  PIN addr_rd_out[55] 
    ANTENNAPARTIALMETALAREA 0.1022 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4088 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.1372 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6272 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal4 ; 
    ANTENNAMAXAREACAR 11.0048 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 41.3657 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.24998 LAYER via4 ;
  END addr_rd_out[55]
  PIN addr_rd_out[54] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2702 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0808 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.5996 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 40.6558 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[54]
  PIN addr_rd_out[53] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3766 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.526 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.72504 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 34.426 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[53]
  PIN addr_rd_out[52] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1841 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7364 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.735 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 52.6156 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[52]
  PIN addr_rd_out[51] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.02695 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1078 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.4513 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.6649 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[51]
  PIN addr_rd_out[50] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.378 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.19349 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.579 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[50]
  PIN addr_rd_out[49] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3269 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3272 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5354 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.1337 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_rd_out[49]
  PIN addr_rd_out[48] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4032 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6324 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.5447 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 58.0644 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_rd_out[48]
  PIN addr_rd_out[47] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.19845 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8134 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.74139 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 33.5659 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[47]
  PIN addr_rd_out[46] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1043 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4172 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.3487 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 40.0598 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[46]
  PIN addr_rd_out[45] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4312 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.63945 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 38.4743 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[45]
  PIN addr_rd_out[44] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0546 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2184 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.4982 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 34.6386 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[44]
  PIN addr_rd_out[43] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2072 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8484 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.7322 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.3933 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_rd_out[43]
  PIN addr_rd_out[42] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1841 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.756 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.5717 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 45.5942 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_rd_out[42]
  PIN addr_rd_out[41] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.14665 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6062 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.27161 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 37.003 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_rd_out[41]
  PIN addr_rd_out[40] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.26285 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0906 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.68806 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 22.6886 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_rd_out[40]
  PIN addr_rd_out[39] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0511 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2044 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.04804 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.9838 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[39]
  PIN addr_rd_out[38] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2107 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 23.832 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 94.2719 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_rd_out[38]
  PIN addr_rd_out[37] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.14945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6174 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.21046 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 32.7584 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_rd_out[37]
  PIN addr_rd_out[36] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1442 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5964 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 3.74926 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 14.9892 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[36]
  PIN addr_rd_out[35] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.02695 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1078 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.51719 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 36.5443 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[35]
  PIN addr_rd_out[34] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1974 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8092 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.6832 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 45.8221 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[34]
  PIN addr_rd_out[33] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2772 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1284 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.379 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 48.3337 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[33]
  PIN addr_rd_out[32] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2471 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0276 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.94572 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 27.8865 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[32]
  PIN addr_rd_out[31] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3332 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.372 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.0639 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 51.9063 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.37512 LAYER via3 ;
  END addr_rd_out[31]
  PIN addr_rd_out[30] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1806 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.742 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 4.52214 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 17.9 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[30]
  PIN addr_rd_out[29] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2205 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9016 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.27558 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 37.1241 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[29]
  PIN addr_rd_out[28] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4865 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9852 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.48723 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 26.0332 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[28]
  PIN addr_rd_out[27] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.7742 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1164 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.4429 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 29.7934 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[27]
  PIN addr_rd_out[26] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3668 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5064 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.8437 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.5214 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_rd_out[26]
  PIN addr_rd_out[25] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4697 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8984 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.2348 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 56.2582 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.37512 LAYER via3 ;
  END addr_rd_out[25]
  PIN addr_rd_out[24] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.329 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.0502 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 50.074 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[24]
  PIN addr_rd_out[23] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.672 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.688 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.452 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 48.3767 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[23]
  PIN addr_rd_out[22] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5033 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0328 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.5646 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 53.4205 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_rd_out[22]
  PIN addr_rd_out[21] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5425 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1896 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.19295 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.6883 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[21]
  PIN addr_rd_out[20] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.7651 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.08 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.3281 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 57.2913 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[20]
  PIN addr_rd_out[19] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1876 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7504 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.29608 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 35.8574 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[19]
  PIN addr_rd_out[18] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.94605 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8038 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.1856 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 40.702 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[18]
  PIN addr_rd_out[17] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8351 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.36 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.8719 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 55.4662 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[17]
  PIN addr_rd_out[16] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8288 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3544 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.43339 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 33.7749 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[16]
  PIN addr_rd_out[15] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4312 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7056 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal4 ; 
    ANTENNAMAXAREACAR 12.0156 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 47.5465 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via4 ;
  END addr_rd_out[15]
  PIN addr_rd_out[14] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.0577 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2308 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.4641 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 52.4251 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[14]
  PIN addr_rd_out[13] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.161 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6636 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 19.8413 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 79.2507 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_rd_out[13]
  PIN addr_rd_out[12] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.00735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0294 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.24055 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 35.8741 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[12]
  PIN addr_rd_out[11] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1211 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4844 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.90983 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.5558 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[11]
  PIN addr_rd_out[10] 
    ANTENNAPARTIALMETALAREA 0.5971 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3884 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal4 ; 
    ANTENNAMAXAREACAR 9.77543 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 39.5176 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via4 ;
  END addr_rd_out[10]
  PIN addr_rd_out[9] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.15885 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6746 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.453 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 53.4626 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_rd_out[9]
  PIN addr_rd_out[8] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.42385 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.715 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.42092 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 25.6625 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[8]
  PIN addr_rd_out[7] 
    ANTENNAPARTIALMETALAREA 0.1106 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4424 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal4 ; 
    ANTENNAMAXAREACAR 12.3371 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 49.9513 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via4 ;
  END addr_rd_out[7]
  PIN addr_rd_out[6] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.43815 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7722 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.7316 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 50.673 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_rd_out[6]
  PIN addr_rd_out[5] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.4805 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9416 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.4543 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 57.7959 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[5]
  PIN addr_rd_out[4] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.25125 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0246 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.5616 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 42.2253 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_rd_out[4]
  PIN addr_rd_out[3] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.11265 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4898 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.5798 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 69.6175 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.37512 LAYER via3 ;
  END addr_rd_out[3]
  PIN addr_rd_out[2] 
    ANTENNAPARTIALMETALAREA 0.0273 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1092 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal4 ; 
    ANTENNAMAXAREACAR 16.0955 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 64.8409 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via4 ;
  END addr_rd_out[2]
  PIN addr_rd_out[1] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3146 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2584 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.1761 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 56.6208 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_rd_out[1]
  PIN addr_rd_out[0] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3811 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5636 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1625 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.6627 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 70.4072 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.169697 LAYER via3 ;
  END addr_rd_out[0]
  PIN addr_wr_out[63] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.15855 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6538 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.13075 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.28695 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 29.0994 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.199793 LAYER via3 ;
  END addr_wr_out[63]
  PIN addr_wr_out[62] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0196 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.10284 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 20.246 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[62]
  PIN addr_wr_out[61] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0196 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.69456 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 26.6129 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[61]
  PIN addr_wr_out[60] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0196 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.64996 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 26.3915 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[60]
  PIN addr_wr_out[59] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1575 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6692 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.0683 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 55.8509 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.37512 LAYER via3 ;
  END addr_wr_out[59]
  PIN addr_wr_out[58] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.18515 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7602 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.03244 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.0463 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[58]
  PIN addr_wr_out[57] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3738 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5148 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.0833 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 47.7862 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_wr_out[57]
  PIN addr_wr_out[56] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.11865 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4942 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.0361 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 67.609 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.37512 LAYER via3 ;
  END addr_wr_out[56]
  PIN addr_wr_out[55] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.21175 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8666 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.41985 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 25.6582 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[55]
  PIN addr_wr_out[54] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.063 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.95443 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.6523 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[54]
  PIN addr_wr_out[53] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1708 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7028 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.57115 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 37.5195 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[53]
  PIN addr_wr_out[52] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2674 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0892 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.67991 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 30.6791 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[52]
  PIN addr_wr_out[51] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.00735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0294 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.38148 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 21.3176 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[51]
  PIN addr_wr_out[50] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.063 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.64372 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 25.4332 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_wr_out[50]
  PIN addr_wr_out[49] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.22505 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9198 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.97664 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.8853 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[49]
  PIN addr_wr_out[48] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.16975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6986 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.86111 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 34.9683 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[48]
  PIN addr_wr_out[47] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.13685 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.567 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.33673 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 32.8727 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[47]
  PIN addr_wr_out[46] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.00735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0294 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.54296 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 26.0065 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[46]
  PIN addr_wr_out[45] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1708 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7028 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.90368 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.5446 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[45]
  PIN addr_wr_out[44] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2569 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0472 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.48244 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 33.8463 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[44]
  PIN addr_wr_out[43] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.13195 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5474 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.49308 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 33.3527 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[43]
  PIN addr_wr_out[42] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.06895 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2758 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.45752 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 28.5444 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[42]
  PIN addr_wr_out[41] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.15855 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6538 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.08147 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 36.3047 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[41]
  PIN addr_wr_out[40] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.00735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0294 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 4.96172 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 18.7794 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[40]
  PIN addr_wr_out[39] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.14525 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6006 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 18.3711 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 72.9374 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_wr_out[39]
  PIN addr_wr_out[38] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.25165 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0262 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.91661 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 26.485 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_wr_out[38]
  PIN addr_wr_out[37] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.31465 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2978 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.07495 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 19.9505 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[37]
  PIN addr_wr_out[36] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.29295 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.211 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.84421 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 31.4938 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[36]
  PIN addr_wr_out[35] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.063 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.65719 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 26.4338 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[35]
  PIN addr_wr_out[34] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.25165 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0262 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.8024 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 50.72 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_wr_out[34]
  PIN addr_wr_out[33] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.063 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.89647 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.4205 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[33]
  PIN addr_wr_out[32] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.08365 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3542 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.78042 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 26.9331 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[32]
  PIN addr_wr_out[31] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23835 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.973 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.70761 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 34.7899 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[31]
  PIN addr_wr_out[30] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.00735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0294 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.42848 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 32.2101 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[30]
  PIN addr_wr_out[29] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09555 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3822 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.79206 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 34.028 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[29]
  PIN addr_wr_out[28] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.19845 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8134 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.18012 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.6503 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[28]
  PIN addr_wr_out[27] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.14525 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6006 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.08744 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 28.2796 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[27]
  PIN addr_wr_out[26] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2205 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9016 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.94647 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 27.7453 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[26]
  PIN addr_wr_out[25] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0196 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.04949 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 31.0084 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_wr_out[25]
  PIN addr_wr_out[24] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1939 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7952 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.51101 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 29.9739 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[24]
  PIN addr_wr_out[23] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1274 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.05921 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.3211 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[23]
  PIN addr_wr_out[22] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.161 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6636 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.96772 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 32.0368 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[22]
  PIN addr_wr_out[21] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.224 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9156 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.65546 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 37.6385 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[21]
  PIN addr_wr_out[20] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0196 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.15783 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.6599 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_wr_out[20]
  PIN addr_wr_out[19] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0196 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.5231 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 21.6921 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[19]
  PIN addr_wr_out[18] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1477 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6104 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.23628 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 28.9046 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[18]
  PIN addr_wr_out[17] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.00735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0294 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.06016 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 28.0753 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[17]
  PIN addr_wr_out[16] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.00735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0294 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.53636 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 28.8391 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_wr_out[16]
  PIN addr_wr_out[15] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.00735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0294 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.90984 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.5988 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[15]
  PIN addr_wr_out[14] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0196 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.16819 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 27.4258 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_wr_out[14]
  PIN addr_wr_out[13] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1841 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.756 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.99328 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 27.9326 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[13]
  PIN addr_wr_out[12] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1309 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5432 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.24647 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.9453 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.1562 LAYER via3 ;
  END addr_wr_out[12]
  PIN addr_wr_out[11] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.01715 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0686 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.09501 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.2919 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[11]
  PIN addr_wr_out[10] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.112 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.07927 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.2765 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[10]
  PIN addr_wr_out[9] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0413 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1652 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.20188 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.6422 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[9]
  PIN addr_wr_out[8] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.112 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.50284 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 25.846 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[8]
  PIN addr_wr_out[7] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.112 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.21096 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 27.5222 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.21877 LAYER via3 ;
  END addr_wr_out[7]
  PIN addr_wr_out[6] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.00735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0294 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.38871 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 21.3599 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[6]
  PIN addr_wr_out[5] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.063 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.07184 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 28.0924 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.12499 LAYER via3 ;
  END addr_wr_out[5]
  PIN addr_wr_out[4] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.14525 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6006 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.63327 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 38.5252 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[4]
  PIN addr_wr_out[3] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.30415 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2558 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.5955 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 34.4856 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[3]
  PIN addr_wr_out[2] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.39445 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.077 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 55.5223 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END addr_wr_out[2]
  PIN addr_wr_out[1] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3976 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.157 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.2284 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 29.0929 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END addr_wr_out[1]
  PIN addr_wr_out[0] 
    ANTENNAPARTIALMETALAREA 0.0567 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2464 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.10475 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.50955 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 30.2635 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.187112 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal4 ;
    ANTENNAGATEAREA 0.10475 LAYER metal4 ; 
    ANTENNAMAXAREACAR 8.44511 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 34.7542 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.374224 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.862 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5264 LAYER metal5 ;
    ANTENNAGATEAREA 0.10475 LAYER metal5 ; 
    ANTENNAMAXAREACAR 26.2208 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 106.605 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 0.561337 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 36.9656 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 148.019 LAYER metal6 ;
    ANTENNAGATEAREA 0.131 LAYER metal6 ; 
    ANTENNAMAXAREACAR 354.38 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1422.66 LAYER metal6 ;
    ANTENNAMAXCUTCAR 2.05333 LAYER via6 ;
  END addr_wr_out[0]
  PIN n_out[127] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 186.25 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 747.651 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.687719 LAYER via7 ;
  END n_out[127]
  PIN n_out[126] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 256.22 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1028.75 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.797129 LAYER via7 ;
  END n_out[126]
  PIN n_out[125] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 568.288 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 2278.65 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[125]
  PIN n_out[124] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 267.537 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1074.24 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.797129 LAYER via7 ;
  END n_out[124]
  PIN n_out[123] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 252.382 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1014.42 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.890909 LAYER via7 ;
  END n_out[123]
  PIN n_out[122] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 519.11 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 2081.56 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[122]
  PIN n_out[121] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 776.341 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 3110.49 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.62552 LAYER via7 ;
  END n_out[121]
  PIN n_out[120] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 247.669 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 997.058 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.21914 LAYER via7 ;
  END n_out[120]
  PIN n_out[119] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 617.594 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 2475.13 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[119]
  PIN n_out[118] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 828.601 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 3318.78 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[118]
  PIN n_out[117] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 408.733 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1639.82 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.59426 LAYER via7 ;
  END n_out[117]
  PIN n_out[116] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 197.57 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 792.57 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.797129 LAYER via7 ;
  END n_out[116]
  PIN n_out[115] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 249.119 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 998.17 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.797129 LAYER via7 ;
  END n_out[115]
  PIN n_out[114] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 379.266 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1523.45 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.59426 LAYER via7 ;
  END n_out[114]
  PIN n_out[113] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 388.544 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1559.06 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.59426 LAYER via7 ;
  END n_out[113]
  PIN n_out[112] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 572.794 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 2295.49 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[112]
  PIN n_out[111] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 358.723 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1439.64 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.30301 LAYER via7 ;
  END n_out[111]
  PIN n_out[110] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 165.692 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 665.472 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.890909 LAYER via7 ;
  END n_out[110]
  PIN n_out[109] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 284.906 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1144.65 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.59426 LAYER via7 ;
  END n_out[109]
  PIN n_out[108] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 212.352 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 854.636 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.30301 LAYER via7 ;
  END n_out[108]
  PIN n_out[107] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[107]
  PIN n_out[106] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 159.121 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 640.76 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.21914 LAYER via7 ;
  END n_out[106]
  PIN n_out[105] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 230.355 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 926.718 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.30301 LAYER via7 ;
  END n_out[105]
  PIN n_out[104] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 270.508 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1092.58 LAYER metal7 ;
    ANTENNAMAXCUTCAR 3.04968 LAYER via7 ;
  END n_out[104]
  PIN n_out[103] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 440.583 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1770.88 LAYER metal7 ;
    ANTENNAMAXCUTCAR 3.04968 LAYER via7 ;
  END n_out[103]
  PIN n_out[102] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 198.909 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 801.012 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[102]
  PIN n_out[101] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 557.451 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 2237.91 LAYER metal7 ;
    ANTENNAMAXCUTCAR 3.04968 LAYER via7 ;
  END n_out[101]
  PIN n_out[100] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 215.868 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 869.11 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.21914 LAYER via7 ;
  END n_out[100]
  PIN n_out[99] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[99]
  PIN n_out[98] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 209.789 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 842.088 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.750239 LAYER via7 ;
  END n_out[98]
  PIN n_out[97] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 244.156 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 982.262 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.59426 LAYER via7 ;
  END n_out[97]
  PIN n_out[96] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 228.89 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 918.76 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.797129 LAYER via7 ;
  END n_out[96]
  PIN n_out[95] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 233.525 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 936.93 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.797129 LAYER via7 ;
  END n_out[95]
  PIN n_out[94] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 236.134 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 947.673 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.750239 LAYER via7 ;
  END n_out[94]
  PIN n_out[93] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 484.869 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1944.08 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.30301 LAYER via7 ;
  END n_out[93]
  PIN n_out[92] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 923.998 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 3705.54 LAYER metal7 ;
    ANTENNAMAXCUTCAR 3.04968 LAYER via7 ;
  END n_out[92]
  PIN n_out[91] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 627.549 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 2518.58 LAYER metal7 ;
    ANTENNAMAXCUTCAR 3.04968 LAYER via7 ;
  END n_out[91]
  PIN n_out[90] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 316.114 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1274.86 LAYER metal7 ;
    ANTENNAMAXCUTCAR 3.04968 LAYER via7 ;
  END n_out[90]
  PIN n_out[89] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 281.77 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1134.45 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.30301 LAYER via7 ;
  END n_out[89]
  PIN n_out[88] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 198.633 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 798.48 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.797129 LAYER via7 ;
  END n_out[88]
  PIN n_out[87] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ; 
    ANTENNAMAXAREACAR 566.788 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 2276.26 LAYER metal7 ;
    ANTENNAMAXCUTCAR 3.04968 LAYER via7 ;
  END n_out[87]
  PIN n_out[86] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 243.107 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 977.035 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.797129 LAYER via7 ;
  END n_out[86]
  PIN n_out[85] 
    ANTENNADIFFAREA 2.3617 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 270.836 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1090.11 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.59426 LAYER via7 ;
  END n_out[85]
  PIN n_out[84] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ; 
    ANTENNAMAXAREACAR 232.099 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 934.783 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.59426 LAYER via7 ;
  END n_out[84]
  PIN n_out[83] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 198.048 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 795.367 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.2504 LAYER via7 ;
  END n_out[83]
  PIN n_out[82] 
    ANTENNADIFFAREA 0.1463 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 409.177 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1642.1 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[82]
  PIN n_out[81] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 182.42 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 735.429 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.2504 LAYER via7 ;
  END n_out[81]
  PIN n_out[80] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 280.723 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1125.47 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[80]
  PIN n_out[79] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 387.474 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1555.45 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[79]
  PIN n_out[78] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 317.655 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1274.78 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[78]
  PIN n_out[77] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 280.67 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1126.98 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[77]
  PIN n_out[76] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 173.759 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 696.908 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.593939 LAYER via7 ;
  END n_out[76]
  PIN n_out[75] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 160.873 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 645.99 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.687719 LAYER via7 ;
  END n_out[75]
  PIN n_out[74] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 196.795 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 791.659 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[74]
  PIN n_out[73] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 173.083 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 694.795 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[73]
  PIN n_out[72] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 164.235 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 658.326 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.687719 LAYER via7 ;
  END n_out[72]
  PIN n_out[71] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 242.345 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 974.63 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.2504 LAYER via7 ;
  END n_out[71]
  PIN n_out[70] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 174.952 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 702.792 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[70]
  PIN n_out[69] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 230.109 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 925.613 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[69]
  PIN n_out[68] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 208.477 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 839.159 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[68]
  PIN n_out[67] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 193.593 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 776.444 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[67]
  PIN n_out[66] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 178.685 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 716.683 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[66]
  PIN n_out[65] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 209.164 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 839.747 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[65]
  PIN n_out[64] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 215.367 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 864.667 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[64]
  PIN n_out[63] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 182.746 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 734.683 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.09442 LAYER via7 ;
  END n_out[63]
  PIN n_out[62] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 205.838 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 827.363 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[62]
  PIN n_out[61] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 199.782 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 803.859 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[61]
  PIN n_out[60] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 218.125 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 877.376 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[60]
  PIN n_out[59] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 218.03 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 874.822 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[59]
  PIN n_out[58] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 206.315 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 828.08 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[58]
  PIN n_out[57] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 231.77 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 935.207 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.09442 LAYER via7 ;
  END n_out[57]
  PIN n_out[56] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 208.857 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 840.802 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[56]
  PIN n_out[55] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 219.941 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 884.064 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[55]
  PIN n_out[54] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 198.9 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 798.174 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.00064 LAYER via7 ;
  END n_out[54]
  PIN n_out[53] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 229.156 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 921.011 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.09442 LAYER via7 ;
  END n_out[53]
  PIN n_out[52] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 281.152 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1129.21 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.53174 LAYER via7 ;
  END n_out[52]
  PIN n_out[51] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 225.695 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 905.356 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.00064 LAYER via7 ;
  END n_out[51]
  PIN n_out[50] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 312.381 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1254.77 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.2504 LAYER via7 ;
  END n_out[50]
  PIN n_out[49] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 262.448 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1054.68 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[49]
  PIN n_out[48] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 218.262 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 874.92 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[48]
  PIN n_out[47] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 234.968 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 942.759 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.15662 LAYER via7 ;
  END n_out[47]
  PIN n_out[46] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ; 
    ANTENNAMAXAREACAR 244.188 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 981.029 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.2504 LAYER via7 ;
  END n_out[46]
  PIN n_out[45] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[45]
  PIN n_out[44] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[44]
  PIN n_out[43] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[43]
  PIN n_out[42] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[42]
  PIN n_out[41] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1081.83 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4339 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[41]
  PIN n_out[40] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[40]
  PIN n_out[39] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[39]
  PIN n_out[38] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[38]
  PIN n_out[37] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[37]
  PIN n_out[36] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[36]
  PIN n_out[35] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1092.24 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4381.48 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[35]
  PIN n_out[34] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[34]
  PIN n_out[33] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[33]
  PIN n_out[32] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[32]
  PIN n_out[31] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[31]
  PIN n_out[30] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1150.2 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4619.15 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[30]
  PIN n_out[29] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1168.73 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4693.43 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[29]
  PIN n_out[28] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1187.37 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4762.76 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[28]
  PIN n_out[27] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1143.33 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4584.99 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[27]
  PIN n_out[26] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1185.23 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4756.42 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[26]
  PIN n_out[25] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ; 
    ANTENNAMAXAREACAR 609.717 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 2446.74 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.4067 LAYER via7 ;
  END n_out[25]
  PIN n_out[24] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1169.17 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4691.91 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[24]
  PIN n_out[23] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1173.05 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4709.07 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[23]
  PIN n_out[22] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1175.29 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4716.68 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[22]
  PIN n_out[21] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1177.05 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4726.71 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[21]
  PIN n_out[20] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[20]
  PIN n_out[19] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[19]
  PIN n_out[18] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1146.99 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4600.5 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[18]
  PIN n_out[17] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1135.67 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4557.74 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[17]
  PIN n_out[16] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[16]
  PIN n_out[15] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1289.48 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 5169.86 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[15]
  PIN n_out[14] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[14]
  PIN n_out[13] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1256.6 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 5041.91 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[13]
  PIN n_out[12] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1241.96 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4983.2 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[12]
  PIN n_out[11] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1221.83 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4899.33 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[11]
  PIN n_out[10] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[10]
  PIN n_out[9] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[9]
  PIN n_out[8] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1232.35 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4941.33 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[8]
  PIN n_out[7] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ; 
    ANTENNAMAXAREACAR 1174.12 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 4709.6 LAYER metal7 ;
    ANTENNAMAXCUTCAR 2.8 LAYER via7 ;
  END n_out[7]
  PIN n_out[6] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
  END n_out[6]
  PIN n_out[5] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.13075 LAYER metal7 ; 
    ANTENNAMAXAREACAR 230.128 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 923.311 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.618445 LAYER via7 ;
  END n_out[5]
  PIN n_out[4] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.183 LAYER metal7 ; 
    ANTENNAMAXAREACAR 203.779 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 818.275 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.870667 LAYER via7 ;
  END n_out[4]
  PIN n_out[3] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.183 LAYER metal7 ; 
    ANTENNAMAXAREACAR 296.579 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 1190.9 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.5138 LAYER via7 ;
  END n_out[3]
  PIN n_out[2] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.183 LAYER metal7 ; 
    ANTENNAMAXAREACAR 193.709 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 777.191 LAYER metal7 ;
    ANTENNAMAXCUTCAR 1.13868 LAYER via7 ;
  END n_out[2]
  PIN n_out[1] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.13075 LAYER metal7 ; 
    ANTENNAMAXAREACAR 230.072 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 922.419 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.618445 LAYER via7 ;
  END n_out[1]
  PIN n_out[0] 
    ANTENNADIFFAREA 0.109725 LAYER metal7 ; 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.13075 LAYER metal7 ; 
    ANTENNAMAXAREACAR 218.954 LAYER metal7 ;
    ANTENNAMAXSIDEAREACAR 878.015 LAYER metal7 ;
    ANTENNAMAXCUTCAR 0.674749 LAYER via7 ;
  END n_out[0]
  PIN g_out[127] 
    ANTENNADIFFAREA 0.1463 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.33565 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3426 LAYER metal3 ;
  END g_out[127]
  PIN g_out[126] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.27265 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0906 LAYER metal3 ;
  END g_out[126]
  PIN g_out[125] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.36575 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER metal3 ;
  END g_out[125]
  PIN g_out[124] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[124]
  PIN g_out[123] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[123]
  PIN g_out[122] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[122]
  PIN g_out[121] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[121]
  PIN g_out[120] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.24605 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9842 LAYER metal3 ;
  END g_out[120]
  PIN g_out[119] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.25935 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0374 LAYER metal3 ;
  END g_out[119]
  PIN g_out[118] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.27545 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1018 LAYER metal3 ;
  END g_out[118]
  PIN g_out[117] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.24255 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9702 LAYER metal3 ;
  END g_out[117]
  PIN g_out[116] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.20615 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8246 LAYER metal3 ;
  END g_out[116]
  PIN g_out[115] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5054 LAYER metal3 ;
  END g_out[115]
  PIN g_out[114] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.21945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8778 LAYER metal3 ;
  END g_out[114]
  PIN g_out[113] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[113]
  PIN g_out[112] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[112]
  PIN g_out[111] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[111]
  PIN g_out[110] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.25235 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0094 LAYER metal3 ;
  END g_out[110]
  PIN g_out[109] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.07315 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER metal3 ;
  END g_out[109]
  PIN g_out[108] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.29225 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.169 LAYER metal3 ;
  END g_out[108]
  PIN g_out[107] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.07315 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER metal3 ;
  END g_out[107]
  PIN g_out[106] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[106]
  PIN g_out[105] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[105]
  PIN g_out[104] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[104]
  PIN g_out[103] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.24605 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9842 LAYER metal3 ;
  END g_out[103]
  PIN g_out[102] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.26565 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0626 LAYER metal3 ;
  END g_out[102]
  PIN g_out[101] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.59815 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3926 LAYER metal3 ;
  END g_out[101]
  PIN g_out[100] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[100]
  PIN g_out[99] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.27265 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0906 LAYER metal3 ;
  END g_out[99]
  PIN g_out[98] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5054 LAYER metal3 ;
  END g_out[98]
  PIN g_out[97] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.08295 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3318 LAYER metal3 ;
  END g_out[97]
  PIN g_out[96] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[96]
  PIN g_out[95] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.27265 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0906 LAYER metal3 ;
  END g_out[95]
  PIN g_out[94] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[94]
  PIN g_out[93] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.60795 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4318 LAYER metal3 ;
  END g_out[93]
  PIN g_out[92] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[92]
  PIN g_out[91] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[91]
  PIN g_out[90] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[90]
  PIN g_out[89] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[89]
  PIN g_out[88] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.47845 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9334 LAYER metal3 ;
  END g_out[88]
  PIN g_out[87] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5054 LAYER metal3 ;
  END g_out[87]
  PIN g_out[86] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.84735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3894 LAYER metal3 ;
  END g_out[86]
  PIN g_out[85] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.60165 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4066 LAYER metal3 ;
  END g_out[85]
  PIN g_out[84] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.22575 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.903 LAYER metal3 ;
  END g_out[84]
  PIN g_out[83] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.27895 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1158 LAYER metal3 ;
  END g_out[83]
  PIN g_out[82] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3458 LAYER metal3 ;
  END g_out[82]
  PIN g_out[81] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[81]
  PIN g_out[80] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[80]
  PIN g_out[79] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.21945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8778 LAYER metal3 ;
  END g_out[79]
  PIN g_out[78] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.31535 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2614 LAYER metal3 ;
  END g_out[78]
  PIN g_out[77] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.02625 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.105 LAYER metal3 ;
  END g_out[77]
  PIN g_out[76] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.28245 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1298 LAYER metal3 ;
  END g_out[76]
  PIN g_out[75] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[75]
  PIN g_out[74] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4522 LAYER metal3 ;
  END g_out[74]
  PIN g_out[73] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[73]
  PIN g_out[72] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[72]
  PIN g_out[71] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.07315 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2926 LAYER metal3 ;
  END g_out[71]
  PIN g_out[70] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.29225 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.169 LAYER metal3 ;
  END g_out[70]
  PIN g_out[69] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[69]
  PIN g_out[68] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.33625 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.345 LAYER metal3 ;
  END g_out[68]
  PIN g_out[67] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.85815 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4326 LAYER metal3 ;
  END g_out[67]
  PIN g_out[66] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.99745 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9898 LAYER metal3 ;
  END g_out[66]
  PIN g_out[65] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.54525 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.181 LAYER metal3 ;
  END g_out[65]
  PIN g_out[64] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.79025 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1806 LAYER metal3 ;
  END g_out[64]
  PIN g_out[63] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.10035 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4014 LAYER metal3 ;
  END g_out[63]
  PIN g_out[62] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.39545 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5818 LAYER metal3 ;
  END g_out[62]
  PIN g_out[61] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.72795 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9314 LAYER metal3 ;
  END g_out[61]
  PIN g_out[60] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.93055 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.7222 LAYER metal3 ;
  END g_out[60]
  PIN g_out[59] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.98315 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9326 LAYER metal3 ;
  END g_out[59]
  PIN g_out[58] 
    ANTENNAPARTIALMETALAREA 1.86585 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4634 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 0.2548 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0976 LAYER metal5 ;
  END g_out[58]
  PIN g_out[57] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.93125 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.725 LAYER metal3 ;
  END g_out[57]
  PIN g_out[56] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 3.26305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0718 LAYER metal3 ;
  END g_out[56]
  PIN g_out[55] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 3.06985 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.299 LAYER metal3 ;
  END g_out[55]
  PIN g_out[54] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.89205 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5682 LAYER metal3 ;
  END g_out[54]
  PIN g_out[53] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.53785 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.171 LAYER metal3 ;
  END g_out[53]
  PIN g_out[52] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.01065 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0622 LAYER metal3 ;
  END g_out[52]
  PIN g_out[51] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.01135 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0454 LAYER metal3 ;
  END g_out[51]
  PIN g_out[50] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.00715 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0286 LAYER metal3 ;
  END g_out[50]
  PIN g_out[49] 
    ANTENNAPARTIALMETALAREA 0.12145 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4858 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 2.0972 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4672 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 0.5292 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1952 LAYER metal6 ;
  END g_out[49]
  PIN g_out[48] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.49795 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9918 LAYER metal3 ;
  END g_out[48]
  PIN g_out[47] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.71565 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8626 LAYER metal3 ;
  END g_out[47]
  PIN g_out[46] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.93125 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.7446 LAYER metal3 ;
  END g_out[46]
  PIN g_out[45] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.03035 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1214 LAYER metal3 ;
  END g_out[45]
  PIN g_out[44] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.05415 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2166 LAYER metal3 ;
  END g_out[44]
  PIN g_out[43] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[43]
  PIN g_out[42] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.21945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8778 LAYER metal3 ;
  END g_out[42]
  PIN g_out[41] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.37905 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5162 LAYER metal3 ;
  END g_out[41]
  PIN g_out[40] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[40]
  PIN g_out[39] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.24605 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9842 LAYER metal3 ;
  END g_out[39]
  PIN g_out[38] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.28245 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1494 LAYER metal3 ;
  END g_out[38]
  PIN g_out[37] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.22925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.917 LAYER metal3 ;
  END g_out[37]
  PIN g_out[36] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[36]
  PIN g_out[35] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[35]
  PIN g_out[34] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.39235 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5694 LAYER metal3 ;
  END g_out[34]
  PIN g_out[33] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23905 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9562 LAYER metal3 ;
  END g_out[33]
  PIN g_out[32] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[32]
  PIN g_out[31] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.29225 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1886 LAYER metal3 ;
  END g_out[31]
  PIN g_out[30] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3458 LAYER metal3 ;
  END g_out[30]
  PIN g_out[29] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1386 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5544 LAYER metal3 ;
  END g_out[29]
  PIN g_out[28] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.27545 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1018 LAYER metal3 ;
  END g_out[28]
  PIN g_out[27] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4522 LAYER metal3 ;
  END g_out[27]
  PIN g_out[26] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.24255 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9702 LAYER metal3 ;
  END g_out[26]
  PIN g_out[25] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.21945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8778 LAYER metal3 ;
  END g_out[25]
  PIN g_out[24] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[24]
  PIN g_out[23] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.08645 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3458 LAYER metal3 ;
  END g_out[23]
  PIN g_out[22] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.34895 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4154 LAYER metal3 ;
  END g_out[22]
  PIN g_out[21] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.29575 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2026 LAYER metal3 ;
  END g_out[21]
  PIN g_out[20] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.23275 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER metal3 ;
  END g_out[20]
  PIN g_out[19] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5054 LAYER metal3 ;
  END g_out[19]
  PIN g_out[18] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.25585 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0234 LAYER metal3 ;
  END g_out[18]
  PIN g_out[17] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.30555 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2222 LAYER metal3 ;
  END g_out[17]
  PIN g_out[16] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.21945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8778 LAYER metal3 ;
  END g_out[16]
  PIN g_out[15] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.09975 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.399 LAYER metal3 ;
  END g_out[15]
  PIN g_out[14] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.21945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8778 LAYER metal3 ;
  END g_out[14]
  PIN g_out[13] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.28245 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1298 LAYER metal3 ;
  END g_out[13]
  PIN g_out[12] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.01995 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0798 LAYER metal3 ;
  END g_out[12]
  PIN g_out[11] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.21945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8778 LAYER metal3 ;
  END g_out[11]
  PIN g_out[10] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5054 LAYER metal3 ;
  END g_out[10]
  PIN g_out[9] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4522 LAYER metal3 ;
  END g_out[9]
  PIN g_out[8] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.26915 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0766 LAYER metal3 ;
  END g_out[8]
  PIN g_out[7] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.12635 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5054 LAYER metal3 ;
  END g_out[7]
  PIN g_out[6] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.20615 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8246 LAYER metal3 ;
  END g_out[6]
  PIN g_out[5] 
    ANTENNAPARTIALMETALAREA 0.12145 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4858 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.666 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7424 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.1463 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 0.686 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8224 LAYER metal6 ;
  END g_out[5]
  PIN g_out[4] 
    ANTENNADIFFAREA 0.1463 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.95175 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.8462 LAYER metal3 ;
  END g_out[4]
  PIN g_out[3] 
    ANTENNAPARTIALMETALAREA 0.61145 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4458 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.8428 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4496 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.1463 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.6464 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7424 LAYER metal6 ;
  END g_out[3]
  PIN g_out[2] 
    ANTENNAPARTIALMETALAREA 0.13125 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.7428 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0496 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.1463 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.332 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 13.4848 LAYER metal6 ;
  END g_out[2]
  PIN g_out[1] 
    ANTENNAPARTIALMETALAREA 0.10185 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4074 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.1463 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.4496 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 13.9552 LAYER metal6 ;
  END g_out[1]
  PIN g_out[0] 
    ANTENNAPARTIALMETALAREA 0.112 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.448 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 7.6244 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 30.576 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.038 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 12.2304 LAYER metal6 ;
  END g_out[0]
  PIN lambda_out[127] 
    ANTENNAPARTIALMETALAREA 0.12285 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4914 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.8428 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4496 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 12.7008 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 50.96 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 144.917 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 584.542 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.4067 LAYER via6 ;
  END lambda_out[127]
  PIN lambda_out[126] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.8428 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4496 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 11.074 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 44.3744 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 121.331 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 489.462 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[126]
  PIN lambda_out[125] 
    ANTENNAPARTIALMETALAREA 0.12285 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4914 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6272 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 9.702 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 39.0432 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 129.302 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 522.848 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.4067 LAYER via6 ;
  END lambda_out[125]
  PIN lambda_out[124] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.4116 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 10.4076 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 41.7088 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 112.543 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 454.308 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[124]
  PIN lambda_out[123] 
    ANTENNAPARTIALMETALAREA 0.31885 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2754 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 1.5484 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.272 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 45.9388 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 185.12 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 0.4508 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8816 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 54.5665 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 221.131 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 7.8988 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 31.6736 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 130.153 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 524.228 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[123]
  PIN lambda_out[122] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4522 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 8.526 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.1824 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 104.899 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 421.229 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[122]
  PIN lambda_out[121] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.2586 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.054 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 26.2316 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 105.154 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 26.6067 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 108.155 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 28.4823 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 117.158 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 7.546 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 30.2624 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 100.693 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 406.75 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[121]
  PIN lambda_out[120] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.66745 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6894 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 20.1225 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 80.4995 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.37512 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 20.4976 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 83.5005 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.750239 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 0.3332 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4112 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 26.8746 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 110.509 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.12536 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.9188 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 27.7536 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 93.0833 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 376.094 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.12536 LAYER via6 ;
  END lambda_out[120]
  PIN lambda_out[119] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3744 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.9598 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 55.401 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 14.3349 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 58.4019 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 0.4116 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 22.2124 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 91.4124 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.4092 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 25.7152 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 84.7435 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 343.112 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[119]
  PIN lambda_out[118] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5971 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.408 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.4995 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 50.3713 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 12.8746 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 53.3722 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 14.7502 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 62.3751 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.9388 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.8336 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 71.5809 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 290.448 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[118]
  PIN lambda_out[117] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.55825 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.233 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 16.5388 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 65.9349 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 16.9139 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 68.9359 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 20.29 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 83.9407 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.586 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.4224 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 73.7445 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 298.509 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[117]
  PIN lambda_out[116] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.33845 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3538 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.2744 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.176 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 7.79713 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 33.0622 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 8.17225 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 36.0632 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.4492 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8752 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 52.2287 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 213.053 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[116]
  PIN lambda_out[115] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.76405 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0954 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 19.8211 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 80.0325 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ; 
    ANTENNAMAXAREACAR 20.7589 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 84.534 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via4 ;
  END lambda_out[115]
  PIN lambda_out[114] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.01395 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0558 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 38.6943 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 154.789 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[114]
  PIN lambda_out[113] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.86065 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4426 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 25.2067 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 100.534 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2144 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ; 
    ANTENNAMAXAREACAR 32.7091 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 131.294 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via4 ;
  END lambda_out[113]
  PIN lambda_out[112] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.02305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1314 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 14.211 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 56.6354 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[112]
  PIN lambda_out[111] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.67475 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7186 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 20.7354 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 82.8364 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[111]
  PIN lambda_out[110] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.32195 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3466 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 20.3067 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 81.801 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[110]
  PIN lambda_out[109] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.89695 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.627 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 29.4234 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 117.994 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[109]
  PIN lambda_out[108] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.96065 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9014 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 29.4033 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 118.174 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[108]
  PIN lambda_out[107] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.83365 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3542 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 24.1651 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 96.4995 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.14067 LAYER via3 ;
  END lambda_out[107]
  PIN lambda_out[106] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.29215 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2078 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 27.2196 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 109.265 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[106]
  PIN lambda_out[105] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.6047 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.4384 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 27.578 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 110.207 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[105]
  PIN lambda_out[104] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.32505 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3394 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 25.6522 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 102.691 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[104]
  PIN lambda_out[103] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.30305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2514 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 20.6885 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 83.1407 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[103]
  PIN lambda_out[102] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.21905 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9154 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 20.8359 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 83.7301 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[102]
  PIN lambda_out[101] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.10285 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4506 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.8493 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 55.1885 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[101]
  PIN lambda_out[100] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.58095 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.363 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 16.5287 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 66.5014 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[100]
  PIN lambda_out[99] 
    ANTENNAPARTIALMETALAREA 0.12285 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4914 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.8036 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2928 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.7036 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.8928 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 74.1665 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 300.79 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[99]
  PIN lambda_out[98] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.7828 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.2096 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 7.1736 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 28.8512 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 99.199 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 401.755 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[98]
  PIN lambda_out[97] 
    ANTENNAPARTIALMETALAREA 0.26005 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0402 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.7628 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.1296 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.5464 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 26.3424 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 75.1646 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 305.546 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[97]
  PIN lambda_out[96] 
    ANTENNAPARTIALMETALAREA 0.36785 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4714 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.6452 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.6592 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.1152 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 24.6176 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 70.3684 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 286.362 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[96]
  PIN lambda_out[95] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.7044 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.9188 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 27.7536 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 103.834 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 419.476 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[95]
  PIN lambda_out[94] 
    ANTENNAPARTIALMETALAREA 0.27965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1186 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.9004 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.68 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.2132 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 24.9312 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 91.0402 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 368.299 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[94]
  PIN lambda_out[93] 
    ANTENNAPARTIALMETALAREA 0.36785 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4714 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 6.6444 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 26.656 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.7424 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 27.1264 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 152.573 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 615.181 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[93]
  PIN lambda_out[92] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7056 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 6.6444 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 26.656 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.1936 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 24.9312 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 143.644 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 579.464 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[92]
  PIN lambda_out[91] 
    ANTENNAPARTIALMETALAREA 0.35805 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4322 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.294 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2544 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.4684 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.952 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.3116 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.3248 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 68.2115 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 277.359 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[91]
  PIN lambda_out[90] 
    ANTENNAPARTIALMETALAREA 0.40705 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6282 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 6.8796 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 27.5968 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.3312 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.4816 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 121.231 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 489.811 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[90]
  PIN lambda_out[89] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 6.8796 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 27.5968 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.5664 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.4224 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 68.044 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 276.76 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[89]
  PIN lambda_out[88] 
    ANTENNAPARTIALMETALAREA 0.35805 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4322 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.1744 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 20.8544 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 131.325 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 530.189 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[88]
  PIN lambda_out[87] 
    ANTENNAPARTIALMETALAREA 0.12285 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4914 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.7436 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.0528 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.3708 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.7184 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 52.5904 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 216 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[87]
  PIN lambda_out[86] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4522 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.0356 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 36.2208 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.2336 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0912 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 52.8316 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 216.201 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[86]
  PIN lambda_out[85] 
    ANTENNAPARTIALMETALAREA 0.27965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1186 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 7.0756 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 28.3808 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.724 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 15.0528 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 68.466 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 278.752 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[85]
  PIN lambda_out[84] 
    ANTENNAPARTIALMETALAREA 0.33845 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3538 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 6.9188 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 27.7536 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.3908 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 13.6416 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 59.711 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 242.982 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[84]
  PIN lambda_out[83] 
    ANTENNAPARTIALMETALAREA 0.27965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1186 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.7804 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 39.2 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.0968 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 12.544 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 79.5522 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 323.083 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[83]
  PIN lambda_out[82] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.26995 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1386 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 66.0579 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 264.806 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END lambda_out[82]
  PIN lambda_out[81] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.51145 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.085 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 63.345 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 253.767 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END lambda_out[81]
  PIN lambda_out[80] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.57585 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.3622 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 56.8139 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 227.671 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END lambda_out[80]
  PIN lambda_out[79] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.76485 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0986 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 61.7775 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 247.497 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END lambda_out[79]
  PIN lambda_out[78] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 8.2516 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 33.0848 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ; 
    ANTENNAMAXAREACAR 103.091 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 414.251 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.515789 LAYER via5 ;
  END lambda_out[78]
  PIN lambda_out[77] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 6.13865 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.5938 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 65.1536 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 261.001 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[77]
  PIN lambda_out[76] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 6.34375 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.3946 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 65.9909 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 264.163 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[76]
  PIN lambda_out[75] 
    ANTENNAPARTIALMETALAREA 0.30905 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2362 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7056 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.1164 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 0.7252 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9792 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 88.9167 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 358.247 LAYER metal6 ;
    ANTENNAMAXCUTCAR 0.703349 LAYER via6 ;
  END lambda_out[75]
  PIN lambda_out[74] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 7.17255 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.749 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 72.1469 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 289.148 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END lambda_out[74]
  PIN lambda_out[73] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 9.27955 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.1378 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 105.526 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 422.302 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END lambda_out[73]
  PIN lambda_out[72] 
    ANTENNAPARTIALMETALAREA 0.34825 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.393 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.7644 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 9.2708 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.1616 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ; 
    ANTENNAMAXAREACAR 111.424 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 447.424 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.515789 LAYER via5 ;
  END lambda_out[72]
  PIN lambda_out[71] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 6.9188 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 27.7536 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.1352 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 20.6976 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 132.551 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 538.831 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.96938 LAYER via6 ;
  END lambda_out[71]
  PIN lambda_out[70] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 10.1724 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.768 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.3904 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.7184 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 72.5789 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 295.204 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[70]
  PIN lambda_out[69] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.2708 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.1616 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.8996 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.6768 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 102.347 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 413.527 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[69]
  PIN lambda_out[68] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 11.7404 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 47.04 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.6056 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.5792 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 77.9646 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 316.746 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[68]
  PIN lambda_out[67] 
    ANTENNAPARTIALMETALAREA 0.30905 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2362 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 10.9564 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 43.904 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.5272 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2656 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 90.7856 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 368.031 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[67]
  PIN lambda_out[66] 
    ANTENNAPARTIALMETALAREA 0.31885 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2754 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7056 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.918 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 35.7504 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 7.0364 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 28.224 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 142.278 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 573.248 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.12536 LAYER via6 ;
  END lambda_out[66]
  PIN lambda_out[65] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.5452 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 38.2592 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.4288 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 25.872 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 97.7589 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 395.91 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[65]
  PIN lambda_out[64] 
    ANTENNAPARTIALMETALAREA 0.41685 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6674 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3328 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.5876 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4288 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 7.7812 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 31.36 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 107.184 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 434.373 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[64]
  PIN lambda_out[63] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 13.3868 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 53.6256 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 7.8792 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 31.6736 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 115.664 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 467.544 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[63]
  PIN lambda_out[62] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7056 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.8396 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 35.4368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 7.4872 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 30.1056 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 138.412 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 558.538 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[62]
  PIN lambda_out[61] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.2156 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9408 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 11.1132 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 44.5312 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 8.5652 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.3392 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 92.6478 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 374.425 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[61]
  PIN lambda_out[60] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.8788 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 35.5936 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 7.9772 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 31.9872 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 125.29 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 505.066 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[60]
  PIN lambda_out[59] 
    ANTENNAPARTIALMETALAREA 0.36785 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4714 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7056 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 10.8388 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 43.4336 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 9.212 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.0048 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 110.567 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 446.85 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[59]
  PIN lambda_out[58] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.6828 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 34.8096 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 9.4276 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 37.7888 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 128.164 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 516.792 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[58]
  PIN lambda_out[57] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6272 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.114 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 36.5344 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 8.6632 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 34.8096 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 132.236 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 533.833 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[57]
  PIN lambda_out[56] 
    ANTENNAPARTIALMETALAREA 0.35805 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4322 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.526 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 34.1824 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 10.0156 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.1408 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 178.068 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 716.105 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[56]
  PIN lambda_out[55] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 7.8204 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 31.36 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 10.4664 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 42.0224 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 181.464 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 730.513 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[55]
  PIN lambda_out[54] 
    ANTENNAPARTIALMETALAREA 0.27965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1186 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 11.8188 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 47.3536 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 10.1724 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.768 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 109.039 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 440.295 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[54]
  PIN lambda_out[53] 
    ANTENNAPARTIALMETALAREA 0.27965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1186 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 9.5256 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 38.2592 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 214.361 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 863.962 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.3308 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 25.4016 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 274.943 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1107.04 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via6 ;
  END lambda_out[53]
  PIN lambda_out[52] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.6828 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 34.8096 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.3308 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 25.4016 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 115.262 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 465.187 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[52]
  PIN lambda_out[51] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.2156 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9408 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 11.6032 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 46.5696 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 233.646 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 941.334 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.7232 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0496 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 288.413 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1161.9 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via6 ;
  END lambda_out[51]
  PIN lambda_out[50] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 11.9168 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 47.824 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 241.162 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 971.125 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.782 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.2064 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 296.492 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1193.2 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via6 ;
  END lambda_out[50]
  PIN lambda_out[49] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 12.5832 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 50.4896 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 245.623 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 989.544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.39 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.6384 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 297.202 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1196.61 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via6 ;
  END lambda_out[49]
  PIN lambda_out[48] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.7412 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 39.0432 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.0564 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 24.4608 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 102.367 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 415.095 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.4067 LAYER via6 ;
  END lambda_out[48]
  PIN lambda_out[47] 
    ANTENNAPARTIALMETALAREA 0.31885 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2754 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6272 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 11.3876 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 45.6288 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 227.189 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 912.128 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.37 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 25.5584 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 288.145 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1156.71 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[47]
  PIN lambda_out[46] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 10.3488 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 41.552 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 221.213 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 891.229 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.174 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 24.7744 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 280.295 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1128.3 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via6 ;
  END lambda_out[46]
  PIN lambda_out[45] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 10.6036 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 42.4928 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.37 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 25.5584 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 79.8804 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 323.659 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[45]
  PIN lambda_out[44] 
    ANTENNAPARTIALMETALAREA 0.30905 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2362 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 10.7604 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 43.12 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0392 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 6.8992 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 27.7536 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 122.376 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 494.392 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[44]
  PIN lambda_out[43] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 10.1332 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.6112 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 215.171 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 863.914 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.782 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.2064 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 270.501 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1085.98 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[43]
  PIN lambda_out[42] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 11.7012 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 46.8832 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 232.166 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 931.745 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.8604 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 23.52 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 288.246 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1156.82 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[42]
  PIN lambda_out[41] 
    ANTENNAPARTIALMETALAREA 0.12285 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4914 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.666 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7424 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 5.5272 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2656 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 244.216 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 981.824 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.4067 LAYER via6 ;
  END lambda_out[41]
  PIN lambda_out[40] 
    ANTENNAPARTIALMETALAREA 0.30905 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2362 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.3724 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 10.29 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 41.2384 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 220.282 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 884.503 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.998 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0704 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 268.11 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1076.56 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[40]
  PIN lambda_out[39] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 10.2116 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.9248 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.9196 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 19.7568 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 75.8612 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 307.583 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[39]
  PIN lambda_out[38] 
    ANTENNAPARTIALMETALAREA 0.28945 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1578 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.49 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0384 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 9.3884 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.632 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 195.504 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 785.391 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.4884 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 238.456 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 957.946 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[38]
  PIN lambda_out[37] 
    ANTENNAPARTIALMETALAREA 0.36785 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4714 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 10.0548 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.2976 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 206.463 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 829.977 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.8612 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 15.5232 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 243.412 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 978.524 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[37]
  PIN lambda_out[36] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.114 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 36.5344 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.3316 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.4048 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 73.4431 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 297.606 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[36]
  PIN lambda_out[35] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.8004 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 35.28 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.116 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 16.6208 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 63.2813 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 258.013 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[35]
  PIN lambda_out[34] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.45055 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.8218 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 69.6282 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 278.438 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.14067 LAYER via3 ;
  END lambda_out[34]
  PIN lambda_out[33] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 9.3296 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.4752 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 186.488 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 752.327 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.9004 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 15.68 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 223.812 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 902.375 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.50048 LAYER via6 ;
  END lambda_out[33]
  PIN lambda_out[32] 
    ANTENNAPARTIALMETALAREA 0.27965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1186 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 9.31 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.3184 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ; 
    ANTENNAMAXAREACAR 103.165 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 414.733 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.515789 LAYER via5 ;
  END lambda_out[32]
  PIN lambda_out[31] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.9212 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7632 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.114 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 36.5344 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.0188 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1536 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 41.089 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 168.419 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[31]
  PIN lambda_out[30] 
    ANTENNAPARTIALMETALAREA 0.27965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1186 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 10.0156 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.1408 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 196.79 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 790.536 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.2932 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2512 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 218.735 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 879.064 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[30]
  PIN lambda_out[29] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.49 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0384 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.6068 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5056 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 132.297 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 532.186 LAYER metal6 ;
    ANTENNAMAXCUTCAR 0.703349 LAYER via6 ;
  END lambda_out[29]
  PIN lambda_out[28] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.9396 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.0188 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.1536 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 83.8526 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 337.338 LAYER metal6 ;
    ANTENNAMAXCUTCAR 0.562679 LAYER via6 ;
  END lambda_out[28]
  PIN lambda_out[27] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.40715 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.6874 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 63.7134 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 255.428 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[27]
  PIN lambda_out[26] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.99415 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0158 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 52.4263 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 210.078 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[26]
  PIN lambda_out[25] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 4.5276 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.1888 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ; 
    ANTENNAMAXAREACAR 100.043 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 402.059 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.515789 LAYER via5 ;
  END lambda_out[25]
  PIN lambda_out[24] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.19055 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.7818 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 60.478 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 240.467 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.23445 LAYER via3 ;
  END lambda_out[24]
  PIN lambda_out[23] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.1625 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.7088 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 54.4124 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 218.224 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[23]
  PIN lambda_out[22] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.43585 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.8022 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 58.4349 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 233.791 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END lambda_out[22]
  PIN lambda_out[21] 
    ANTENNAPARTIALMETALAREA 0.27965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1186 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 9.0748 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 36.3776 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 183.916 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 739.122 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.9796 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9968 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 202.859 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 815.646 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[21]
  PIN lambda_out[20] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.91295 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.6518 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 99.0115 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 395.462 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 99.3866 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 398.463 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 3.5084 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.112 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 166.533 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 668.549 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.1756 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.7808 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 187.352 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 752.576 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[20]
  PIN lambda_out[19] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.294 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2544 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.1548 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.6976 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 0.686 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8224 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 42.1876 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 170.938 LAYER metal6 ;
    ANTENNAMAXCUTCAR 0.703349 LAYER via6 ;
  END lambda_out[19]
  PIN lambda_out[18] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 7.40705 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.6674 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 72.9708 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 291.966 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[18]
  PIN lambda_out[17] 
    ANTENNAPARTIALMETALAREA 0.30905 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2362 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 5.1548 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.6976 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 143.068 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 575.646 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.7052 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8992 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 159.386 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 641.667 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[17]
  PIN lambda_out[16] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.0824 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3296 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 81.977 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 327.918 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 82.3522 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 330.919 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 82.7273 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 333.92 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.274 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1744 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 94.9187 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 383.435 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[16]
  PIN lambda_out[15] 
    ANTENNAPARTIALMETALAREA 0.33845 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3538 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.4888 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 14.112 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 127.916 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 516.913 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[15]
  PIN lambda_out[14] 
    ANTENNAPARTIALMETALAREA 0.33845 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3538 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.3328 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4096 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 32.5751 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 132.188 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.3132 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3312 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 57.7081 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 234.22 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.7836 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2128 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 115.282 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 465.108 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[14]
  PIN lambda_out[13] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.32355 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.3334 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 49.8742 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 199.215 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[13]
  PIN lambda_out[12] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.35805 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4322 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 32.0392 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 128.76 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.6076 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5088 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ; 
    ANTENNAMAXAREACAR 37.8536 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 152.767 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via4 ;
  END lambda_out[12]
  PIN lambda_out[11] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.77735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1486 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.4129 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.5885 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[11]
  PIN lambda_out[10] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.92365 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7338 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.2388 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 41.3416 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[10]
  PIN lambda_out[9] 
    ANTENNAPARTIALMETALAREA 0.46865 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8746 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.066 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 44.2756 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 13.3167 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 54.7789 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.234 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0144 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 75.2115 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 303.858 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.7444 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 7.056 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 91.9043 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 371.38 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[9]
  PIN lambda_out[8] 
    ANTENNAPARTIALMETALAREA 0.93625 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7646 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 23.1368 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 92.934 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAMAXCUTCAR 0.37512 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 23.512 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 95.9349 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAMAXCUTCAR 0.750239 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.4292 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7952 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 127.42 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 513.068 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.12536 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.8228 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3696 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 144.863 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 583.59 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.12536 LAYER via6 ;
  END lambda_out[8]
  PIN lambda_out[7] 
    ANTENNAPARTIALMETALAREA 0.32865 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3146 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.7056 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9008 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.5868 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4256 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 71.8689 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 290.863 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.3324 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 9.408 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 94.1885 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 380.892 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[7]
  PIN lambda_out[6] 
    ANTENNAPARTIALMETALAREA 0.29925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6256 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 8.0556 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 32.3008 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 156.967 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 631.633 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 0.6076 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5088 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 162.782 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 655.64 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END lambda_out[6]
  PIN lambda_out[5] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.33855 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.3738 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 61.1144 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 244.425 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[5]
  PIN lambda_out[4] 
    ANTENNAPARTIALMETALAREA 0.37765 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.3524 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.7832 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2896 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 180.433 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 726.532 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.4067 LAYER via6 ;
  END lambda_out[4]
  PIN lambda_out[3] 
    ANTENNAPARTIALMETALAREA 0.41685 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6674 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.4108 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7216 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 65.0531 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 262.431 LAYER metal6 ;
    ANTENNAMAXCUTCAR 0.609569 LAYER via6 ;
  END lambda_out[3]
  PIN lambda_out[2] 
    ANTENNAPARTIALMETALAREA 0.11305 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4522 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.1556 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7008 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 74.0526 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 298.647 LAYER metal6 ;
    ANTENNAMAXCUTCAR 0.609569 LAYER via6 ;
  END lambda_out[2]
  PIN lambda_out[1] 
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.97615 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9438 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.6005 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 42.7751 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END lambda_out[1]
  PIN lambda_out[0] 
    ANTENNAPARTIALMETALAREA 0.27965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1186 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.4492 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8752 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ; 
    ANTENNAMAXAREACAR 96.9952 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 389.981 LAYER metal6 ;
    ANTENNAMAXCUTCAR 0.609569 LAYER via6 ;
  END lambda_out[0]
  PIN u_out[127] 
    ANTENNAPARTIALMETALAREA 0.4137 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5366 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.0395 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1776 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.0763 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3248 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 3.92153 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 15.4756 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[127]
  PIN u_out[126] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4116 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.5725 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3292 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 50.9455 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 203.946 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[126]
  PIN u_out[125] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1764 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8141 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2956 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.8545 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 71.5828 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[125]
  PIN u_out[124] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.5488 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.254 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2093 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8568 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.34258 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 33.1598 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[124]
  PIN u_out[123] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2618 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0668 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.9506 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8416 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 22.3895 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 89.7225 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[123]
  PIN u_out[122] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1764 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.2096 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8776 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 24.4861 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 98.1091 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[122]
  PIN u_out[121] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1736 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.714 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3461 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.404 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 38.312 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 153.037 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[121]
  PIN u_out[120] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.4427 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.81 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 38.9081 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 155.797 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[120]
  PIN u_out[119] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.5519 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2272 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 52.9684 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 212.038 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[119]
  PIN u_out[118] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3332 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.6716 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.706 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 42.1033 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 168.203 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[118]
  PIN u_out[117] 
    ANTENNAPARTIALMETALAREA 0.0546 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2028 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.8694 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4972 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3692 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4964 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 27.7282 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 110.702 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[117]
  PIN u_out[116] 
    ANTENNAPARTIALMETALAREA 0.01715 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2548 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 1.7766 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.126 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6272 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.5876 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4288 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 50.0344 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 204.804 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.12536 LAYER via6 ;
  END u_out[116]
  PIN u_out[115] 
    ANTENNAPARTIALMETALAREA 0.0546 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2028 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.52605 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1238 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.6079 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4904 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 32.1091 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 128.976 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[115]
  PIN u_out[114] 
    ANTENNAPARTIALMETALAREA 0.01715 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1372 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.505 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0788 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 30.3742 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 122.036 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[114]
  PIN u_out[113] 
    ANTENNAPARTIALMETALAREA 0.01715 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.49 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.5484 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2328 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 33.5962 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 134.549 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[113]
  PIN u_out[112] 
    ANTENNAPARTIALMETALAREA 0.0945 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.351 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4116 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.456 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8632 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 30.3943 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 121.742 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[112]
  PIN u_out[111] 
    ANTENNAPARTIALMETALAREA 0.0945 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.351 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2912 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1844 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.1396 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5976 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 26.777 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 107.273 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[111]
  PIN u_out[110] 
    ANTENNAPARTIALMETALAREA 0.0945 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.351 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.8274 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3292 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.12 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4996 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 30.2268 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 120.697 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[110]
  PIN u_out[109] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.12 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5388 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2492 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0164 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 6.29282 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 24.9608 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[109]
  PIN u_out[108] 
    ANTENNAPARTIALMETALAREA 0.2142 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7956 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.147 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6076 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8904 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6008 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 22.1952 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 88.9455 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[108]
  PIN u_out[107] 
    ANTENNAPARTIALMETALAREA 0.0679 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2522 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.294 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1956 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8372 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.388 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.3589 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 69.6 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[107]
  PIN u_out[106] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1225 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5096 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.2761 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1436 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 33.8641 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 135.996 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[106]
  PIN u_out[105] 
    ANTENNAPARTIALMETALAREA 0.2142 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7956 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3598 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3356 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4012 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 27.0852 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 108.88 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[105]
  PIN u_out[104] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1666 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.686 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.7703 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1204 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 36.155 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 144.785 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[104]
  PIN u_out[103] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0882 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3724 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.0468 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2264 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 42.5722 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 170.454 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[103]
  PIN u_out[102] 
    ANTENNAPARTIALMETALAREA 0.0679 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2522 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8036 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.17 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.7192 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 51.5818 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 206.492 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[102]
  PIN u_out[101] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3108 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2628 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.4892 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.996 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 54.2211 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 217.049 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[101]
  PIN u_out[100] 
    ANTENNAPARTIALMETALAREA 0.0546 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2028 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6993 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8168 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.513 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0912 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 49.4316 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 197.891 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[100]
  PIN u_out[99] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.9988 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.0344 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 59.1512 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 236.769 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[99]
  PIN u_out[98] 
    ANTENNAPARTIALMETALAREA 0.01715 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.049 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2156 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.4794 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9568 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 51.6689 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 206.84 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[98]
  PIN u_out[97] 
    ANTENNAPARTIALMETALAREA 0.0945 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.351 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.9964 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0444 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 42.867 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 172.008 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[97]
  PIN u_out[96] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1372 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.9572 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 38.9818 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 156.092 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[96]
  PIN u_out[95] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4116 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.0888 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.3944 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 41.5005 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 166.167 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[95]
  PIN u_out[94] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.147 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6076 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.4882 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0116 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 30.2402 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 121.5 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[94]
  PIN u_out[93] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3332 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.2327 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9896 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 25.1158 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 101.003 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[93]
  PIN u_out[92] 
    ANTENNAPARTIALMETALAREA 0.0679 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2522 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4774 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9292 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.2922 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.208 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 26.6967 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 106.951 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[92]
  PIN u_out[91] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2912 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1844 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8435 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4132 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 22.7445 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 91.1426 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[91]
  PIN u_out[90] 
    ANTENNAPARTIALMETALAREA 0.05565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2067 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.8162 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2844 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.1025 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4296 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 25.1292 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 100.306 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[90]
  PIN u_out[89] 
    ANTENNAPARTIALMETALAREA 0.2142 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7956 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.0556 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2812 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1162 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4844 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 4.87273 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 19.2804 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[89]
  PIN u_out[88] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1372 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8337 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3936 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 18.2967 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 73.7263 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[88]
  PIN u_out[87] 
    ANTENNAPARTIALMETALAREA 0.0945 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.351 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.2558 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0428 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.7609 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0632 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.9081 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 71.422 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[87]
  PIN u_out[86] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3349 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3984 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 26.8842 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 108.077 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[86]
  PIN u_out[85] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5299 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1392 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4487 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8144 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 25.1225 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 100.279 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[85]
  PIN u_out[84] 
    ANTENNAPARTIALMETALAREA 0.06895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2561 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.8288 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3348 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5313 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1644 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.6919 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 46.9321 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[84]
  PIN u_out[83] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.7189 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8952 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5012 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0636 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 11.1627 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 45.1904 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[83]
  PIN u_out[82] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2989 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2152 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8568 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.486 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.9684 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 72.4134 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[82]
  PIN u_out[81] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.12 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4996 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5285 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1336 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 16.5952 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 66.1703 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[81]
  PIN u_out[80] 
    ANTENNAPARTIALMETALAREA 0.05565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2067 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5089 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0552 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.6972 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.828 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 15.4297 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 61.8833 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[80]
  PIN u_out[79] 
    ANTENNAPARTIALMETALAREA 0.05565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2067 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.029 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1356 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3052 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.26 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 10.178 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 40.8766 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[79]
  PIN u_out[78] 
    ANTENNAPARTIALMETALAREA 0.09555 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3549 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.4497 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.838 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.16135 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.40861 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 21.4239 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[78]
  PIN u_out[77] 
    ANTENNAPARTIALMETALAREA 0.09555 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3549 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.64955 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.6178 LAYER metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ; 
    ANTENNAMAXAREACAR 32.7187 LAYER metal2 ;
    ANTENNAMAXSIDEAREACAR 130.289 LAYER metal2 ;
    ANTENNAMAXCUTCAR 0.0937799 LAYER via2 ;
  END u_out[77]
  PIN u_out[76] 
    ANTENNAPARTIALMETALAREA 0.02905 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1079 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.7441 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.996 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1694 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6972 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 23.1129 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 92.2411 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[76]
  PIN u_out[75] 
    ANTENNAPARTIALMETALAREA 0.04235 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1573 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5439 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1952 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.8169 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3264 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 24.9416 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 100.306 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[75]
  PIN u_out[74] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.0668 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2868 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.063 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2716 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 16.9502 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 67.5904 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[74]
  PIN u_out[73] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4501 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.82 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3248 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3384 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.55215 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 30.3732 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[73]
  PIN u_out[72] 
    ANTENNAPARTIALMETALAREA 0.05565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2067 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4823 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9488 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.1722 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.728 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 0.9604 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.92 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 27.5809 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 114.989 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END u_out[72]
  PIN u_out[71] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.0241 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.116 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1526 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6496 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.13301 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 36.6967 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[71]
  PIN u_out[70] 
    ANTENNAPARTIALMETALAREA 0.05565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2067 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.9544 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8372 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8092 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 8.06794 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 32.4364 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via3 ;
  END u_out[70]
  PIN u_out[69] 
    ANTENNAPARTIALMETALAREA 0.09555 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3549 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.3195 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.2976 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2191 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9156 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 5.71675 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 23.0316 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[69]
  PIN u_out[68] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.8778 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5308 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5943 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4164 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 12.8976 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 51.755 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[68]
  PIN u_out[67] 
    ANTENNAPARTIALMETALAREA 0.06895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2561 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4396 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.778 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3657 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5216 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 34.8689 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 140.39 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[67]
  PIN u_out[66] 
    ANTENNAPARTIALMETALAREA 0.09555 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3549 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.9166 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7056 LAYER metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ; 
    ANTENNAMAXAREACAR 37.8297 LAYER metal2 ;
    ANTENNAMAXSIDEAREACAR 151.108 LAYER metal2 ;
    ANTENNAMAXCUTCAR 0.0937799 LAYER via2 ;
  END u_out[66]
  PIN u_out[65] 
    ANTENNAPARTIALMETALAREA 0.06895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2561 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.7469 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0072 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0119 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0672 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5292 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1952 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.0972 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4672 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 57.778 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 235.778 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END u_out[65]
  PIN u_out[64] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1316 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 4.5276 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 18.1888 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 97.3464 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 393.677 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END u_out[64]
  PIN u_out[63] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2541 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2219 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9072 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8624 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5684 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.352 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.8028 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2896 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 83.7282 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 339.204 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END u_out[63]
  PIN u_out[62] 
    ANTENNAPARTIALMETALAREA 0.09555 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3549 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.6884 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7928 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.6041 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4556 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.9885 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 72.1187 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[62]
  PIN u_out[61] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.5813 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3448 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.3752 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5204 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.1923 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 52.5589 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[61]
  PIN u_out[60] 
    ANTENNAPARTIALMETALAREA 0.06895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2561 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6531 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0735 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.2156 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9408 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 22.6641 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 93.0718 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via4 ;
  END u_out[60]
  PIN u_out[59] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6489 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6152 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0588 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.098 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4704 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.4108 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7216 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 64.7445 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 263.644 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END u_out[59]
  PIN u_out[58] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4102 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6604 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.3395 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3776 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.6652 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7392 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 3.5084 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 14.112 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 101.54 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 410.45 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END u_out[58]
  PIN u_out[57] 
    ANTENNAPARTIALMETALAREA 0.06895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2561 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.41645 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.705 LAYER metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ; 
    ANTENNAMAXAREACAR 28.2574 LAYER metal2 ;
    ANTENNAMAXSIDEAREACAR 112.819 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.1162 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4844 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 30.4813 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 122.09 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[57]
  PIN u_out[56] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.3426 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4096 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.2359 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9632 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 7.98086 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 31.7129 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[56]
  PIN u_out[55] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.0353 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1608 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.4021 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6476 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 28.733 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 115.097 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[55]
  PIN u_out[54] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0735 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.9863 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.004 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 21.9005 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 88.1416 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[54]
  PIN u_out[53] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0931 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.917 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7072 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 20.1388 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 80.7196 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[53]
  PIN u_out[52] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3479 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4112 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.6713 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7048 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 1.1956 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8608 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 32.6718 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 131.977 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via4 ;
  END u_out[52]
  PIN u_out[51] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.9891 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.976 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.1361 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5836 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 23.0794 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 92.4823 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[51]
  PIN u_out[50] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.9366 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.766 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.1893 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.816 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 24.2852 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 97.6804 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[50]
  PIN u_out[49] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1715 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7056 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.6086 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4736 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 35.4249 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 141.864 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[49]
  PIN u_out[48] 
    ANTENNAPARTIALMETALAREA 0.02905 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1079 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6685 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6936 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.0272 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.148 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 40.3215 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 161.451 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[48]
  PIN u_out[47] 
    ANTENNAPARTIALMETALAREA 0.05565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2067 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5019 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0272 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.373 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.5312 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 52.3187 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 209.439 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[47]
  PIN u_out[46] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5572 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.268 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.6716 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7452 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 33.5158 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 134.603 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[46]
  PIN u_out[45] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0539 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.6453 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.6204 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 73.0172 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 292.233 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[45]
  PIN u_out[44] 
    ANTENNAPARTIALMETALAREA 0.04235 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1573 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5733 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3128 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.7881 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2112 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 56.9943 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 228.517 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[44]
  PIN u_out[43] 
    ANTENNAPARTIALMETALAREA 0.09555 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3549 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6713 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7244 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 2.8714 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5052 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 65.1665 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 260.456 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[43]
  PIN u_out[42] 
    ANTENNAPARTIALMETALAREA 0.01715 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 1.48785 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0102 LAYER metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ; 
    ANTENNAMAXAREACAR 29.6239 LAYER metal2 ;
    ANTENNAMAXSIDEAREACAR 118.66 LAYER metal2 ;
    ANTENNAMAXCUTCAR 0.0937799 LAYER via2 ;
  END u_out[42]
  PIN u_out[41] 
    ANTENNAPARTIALMETALAREA 0.0945 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.351 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.196 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 3.15245 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7274 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 61.9043 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 249.282 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[41]
  PIN u_out[40] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1176 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.49 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.8029 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2312 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 2.5676 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3488 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 139.293 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 561.837 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.03158 LAYER via6 ;
  END u_out[40]
  PIN u_out[39] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1666 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.686 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 3.9844 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9964 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 77.7799 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 311.659 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[39]
  PIN u_out[38] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5166 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.086 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.5619 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2868 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 91.6459 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 366.748 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[38]
  PIN u_out[37] 
    ANTENNAPARTIALMETALAREA 0.06895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2561 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6461 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.604 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.4828 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 89.489 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 358.496 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[37]
  PIN u_out[36] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2401 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.98 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.7621 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0876 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 93.9234 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 375.858 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[36]
  PIN u_out[35] 
    ANTENNAPARTIALMETALAREA 0.05565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2067 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3087 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2544 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.3164 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2852 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4116 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7248 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 9.2708 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 37.1616 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 189.472 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 761.053 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via5 ;
  END u_out[35]
  PIN u_out[34] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0378 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1708 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.4369 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7672 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 126.566 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 506.052 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[34]
  PIN u_out[33] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.5607 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2624 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 4.9875 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.0284 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 97.0249 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 389.014 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[33]
  PIN u_out[32] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 1.1102 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.48 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.7707 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.122 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 20.6679 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 82.8364 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[32]
  PIN u_out[31] 
    ANTENNAPARTIALMETALAREA 0.5866 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1788 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.7196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.898 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.2052 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.86 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 103.77 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 415.246 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[31]
  PIN u_out[30] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4893 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9768 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 6.2433 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.0516 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 121.83 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 488.233 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[30]
  PIN u_out[29] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2373 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9688 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 6.2881 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.2504 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 121.682 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 488.019 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[29]
  PIN u_out[28] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.525 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1196 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 6.8642 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.4764 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 142.481 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 569.715 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[28]
  PIN u_out[27] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.6069 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4472 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 7.3612 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.5036 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 142.408 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 570.17 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[27]
  PIN u_out[26] 
    ANTENNAPARTIALMETALAREA 0.04235 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1573 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1519 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6272 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.9446 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.8176 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 40.4957 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 162.147 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[26]
  PIN u_out[25] 
    ANTENNAPARTIALMETALAREA 0.09555 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3549 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0637 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2744 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 7.00595 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.063 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 139.849 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 559.935 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[25]
  PIN u_out[24] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1225 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5096 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 8.1053 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.48 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 156.836 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 627.885 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[24]
  PIN u_out[23] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2499 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0192 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 9.4311 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.7832 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 186.076 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 744.842 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[23]
  PIN u_out[22] 
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0931 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.392 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 5.278 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1904 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 102.35 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 410.316 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[22]
  PIN u_out[21] 
    ANTENNAPARTIALMETALAREA 0.06895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2561 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0735 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.3524 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.4684 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 27.4536 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 110.354 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[21]
  PIN u_out[20] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6944 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 10.2466 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.0648 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 197.443 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 790.687 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[20]
  PIN u_out[19] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.42 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6996 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 11.3799 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.5392 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 224.773 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 898.882 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[19]
  PIN u_out[18] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0637 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2744 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.5481 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.212 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 17.8947 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 71.7435 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[18]
  PIN u_out[17] 
    ANTENNAPARTIALMETALAREA 0.05565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2067 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1029 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4312 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 6.8817 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.5464 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 149.294 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 597.34 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[17]
  PIN u_out[16] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2597 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0584 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 11.41 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.6596 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 230.782 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 923.292 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[16]
  PIN u_out[15] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1316 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.3528 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4896 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 263.156 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 1053.91 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via4 ;
  END u_out[15]
  PIN u_out[14] 
    ANTENNAPARTIALMETALAREA 0.09555 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3549 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0735 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3136 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 13.5268 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.1464 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 260.41 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 1041.8 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[14]
  PIN u_out[13] 
    ANTENNAPARTIALMETALAREA 0.0049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0343 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1568 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 8.2642 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.0764 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 174.4 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 697.765 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[13]
  PIN u_out[12] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2891 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.176 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2674 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0892 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6272 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 24.0492 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 96.2752 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 504.492 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 2020.76 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via5 ;
  END u_out[12]
  PIN u_out[11] 
    ANTENNAPARTIALMETALAREA 13.4141 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 49.8238 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.6832 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7524 LAYER metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ; 
    ANTENNAMAXAREACAR 14.2239 LAYER metal2 ;
    ANTENNAMAXSIDEAREACAR 56.31 LAYER metal2 ;
    ANTENNAMAXCUTCAR 0.0937799 LAYER via2 ;
  END u_out[11]
  PIN u_out[10] 
    ANTENNAPARTIALMETALAREA 0.0147 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0546 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.3794 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5568 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 0.4018 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6268 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.02584 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 35.8928 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[10]
  PIN u_out[9] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1568 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6468 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 11.9231 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.7512 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 229.529 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 918.656 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[9]
  PIN u_out[8] 
    ANTENNAPARTIALMETALAREA 0.0413 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1534 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNADIFFAREA 0.109725 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 0.6832 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.772 LAYER metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ; 
    ANTENNAMAXAREACAR 14.2239 LAYER metal2 ;
    ANTENNAMAXSIDEAREACAR 56.6852 LAYER metal2 ;
    ANTENNAMAXCUTCAR 0.0937799 LAYER via2 ;
  END u_out[8]
  PIN u_out[7] 
    ANTENNAPARTIALMETALAREA 0.0413 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1534 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.1274 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 3.4132 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.692 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 82.844 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 331.541 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[7]
  PIN u_out[6] 
    ANTENNAPARTIALMETALAREA 0.08225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.4459 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8032 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 8.4322 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.7484 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNADIFFAREA 0.109725 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 0.6076 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5088 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ; 
    ANTENNAMAXAREACAR 60.8995 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 245.263 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.28134 LAYER via4 ;
  END u_out[6]
  PIN u_out[5] 
    ANTENNAPARTIALMETALAREA 0.1211 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4498 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2646 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.078 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 3.5042 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.0364 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2352 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 3.6652 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7392 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via5 ;
    ANTENNADIFFAREA 0.109725 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1.5876 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4288 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ; 
    ANTENNAMAXAREACAR 266.8 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 1071.87 LAYER metal6 ;
    ANTENNAMAXCUTCAR 1.12536 LAYER via6 ;
  END u_out[5]
  PIN u_out[4] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.2842 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1564 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 11.1251 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.5788 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 214.256 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 857.941 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[4]
  PIN u_out[3] 
    ANTENNAPARTIALMETALAREA 0.0147 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0546 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0784 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3332 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 3.0478 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.25 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 59.667 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 239.208 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[3]
  PIN u_out[2] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 8.4875 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.0284 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 164.714 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 659.77 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[2]
  PIN u_out[1] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0392 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1764 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 3.5903 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3808 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.7836 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.2128 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER via4 ;
    ANTENNADIFFAREA 0.109725 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 9.898 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 39.6704 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ; 
    ANTENNAMAXAREACAR 236.857 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 950.22 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.656459 LAYER via5 ;
  END u_out[1]
  PIN u_out[0] 
    ANTENNAPARTIALMETALAREA 0.1078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4004 LAYER metal1 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER via2 ;
    ANTENNADIFFAREA 0.109725 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 9.8749 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.6172 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ; 
    ANTENNAMAXAREACAR 191.589 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 768.019 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.18756 LAYER via3 ;
  END u_out[0]
END key_generation

END LIBRARY
